<svg width="16" height="13" viewBox="0 0 16 13" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M6.39623 1L1 6.5M1 6.5L6.39623 12M1 6.5H15" stroke="#2CCDA0" stroke-width="1.8" stroke-linecap="round" stroke-linejoin="round"/>
</svg>
